package decoder_pkg;
    /* define enum */
    typedef enum logic[3:0]{
        R, I, S, B, U, J
    } imm_type_t;
    typedef enum logic[8:0]{
        LUI, AUIPC, JAL, JALR, BEQ, BNE, BLT, BGE, BLTU, BGEU,
        LB, LH, LW, LBU, LHU, SB, SH, SW, ADDI, SLTI,
        SLTIU, XORI, ORI, ANDI, ADD, SUB, SLL, SLT, SLTU, XOR,
        SRL, SRA, OR, AND, LWU, LD, SD, SLLI, SRLI, SRAI,
        ADDIW, SLLIW, SRLIW, SRAIW, ADDW, SUBW, SLLW, SRLW, SRAW, FENCE,
        ECALL, EBREAK, MRET, SRET, CSRRW, CSRRS, CSRRC, CSRRWI, CSRRSI, CSRRCI,
        MUL, MULH, MULHSU, MULHU, DIV, DIVU, REM, REMU, MULW, DIVW,
        DIVUW, REMW, REMUW, LRW, SCW, AMOSWAPW, AMOADDW, AMOXORW, AMOANDW, AMOORW,
        AMOMINW, AMOMAXW, AMOMINUW, AMOMAXUW, LRD, SCD, AMOSWAPD, AMOADDD, AMOXORD, AMOANDD,
        AMOORD, AMOMIND, AMOMAXD, AMOMINUD, AMOMAXUD, FLW, FSW, FMADDS, FMSUBS, FNMSUBS,
        FNMADDS, FADDS, FSUBS, FMULS, FDIVS, FSQRTS, FSGNJS, FSGNJNS, FSGNJXS, FMINS,
        FMAXS, FCVTWS, FCVTWUS, FMVXW, FEQS, FLTS, FLES, FCLASSS, FCVTSW, FCVTSWU,
        FMVWX, FCVTLS, FCVTLUS, FCVTSL, FCVTSLU, FLD, FSD, FMADDD, FMSUBD, FNMSUBD,
        FNMADDD, FADDD, FSUBD, FMULD, FDIVD, FSQRTD, FSGNJD, FSGNJND, FSGNJXD, FMIND,
        FMAXD, FCVTSD, FCVTDS, FEQD, FLTD, FLED, FCLASSD, FCVTWD, FCVTWUD, FCVTDW,
        FCVTDWU, FCVTLD, FCVTLUD, FMVXD, FCVTDL, FCVTDLU, FMVDX, FLQ, FSQ, FMADDQ,
        FMSUBQ, FNMSUBQ, FNMADDQ, FADDQ, FSUBQ, FMULQ, FDIVQ, FSQRTQ, FSGNJQ, FSGNJNQ,
        FSGNJXQ, FMINQ, FMAXQ, FCVTSQ, FCVTQS, FCVTDQ, FCVTQD, FEQQ, FLTQ, FLEQ,
        FCLASSQ, FCVTWQ, FCVTWUQ, FCVTQW, FCVTQWU, FCVTLQ, FCVTLUQ, FCVTQL, FCVTQLU, FLH,
        FSH, FMADDH, FMSUBH, FNMSUBH, FNMADDH, FADDH, FSUBH, FMULH, FDIVH, FSQRTH,
        FSGNJH, FSGNJNH, FSGNJXH, FMINH, FMAXH, FCVTSH, FCVTDH, FCVTQH, FCVTHS, FCVTHD,
        FCVTHQ, FMVXH, FEQH, FLTH, FLEH, FCLASSH, FCVTWH, FCVTWUH, FCVTHW, FCVTHWU,
        FMVHX
    } uop_t;
endpackage
